module bfrvlog

pub fn hello() {
	println('hello !')
}
